`define ALU_CTRL_WIDTH 5
`define INSTRUCTION_WIDTH 32

//operand width
`define OPERAND_WIDTH 32
`define IMM_WIDTH 21

`define SIGN_EXTEND 1'b1
`define ZERO_EXTEND 1'b0


//Define the states
//s0 through s23
`define FETCH 0
`define LOAD_IR 1
`define DECODE 2
`define BRANCH_S 3
`define BCOND1 4
`define JALR_S 5
`define JALR2 6
`define JAL_S 7
`define JAL2 8
`define ALU2PC 9
`define AUIPC_S 10
`define WRITE_BACK 11
`define LUI_S 12
`define STORE_S 13
`define STORE_MEM 14
`define LOAD_S 15
`define LOAD2 16
`define I_TYPE_S 17
`define R_TYPE_S 18
`define JALR_ADD 19
`define LOAD_MDR 20
`define LOAD_WR 21
`define PC_ADD 22
`define PC_WR 23

//Define the opcodes for each instruction type
//U-TYPE
`define LUI 5'b01101
`define AUIPC 5'b00101
`define JAL 5'b11011
`define JALR 5'b11001
`define BRANCH 5'b11000
`define LOAD 5'b00000
`define STORE 5'b01000
`define I_TYPE 5'b00100
`define R_TYPE 5'b01100

module cntl_mc_tb;

	// Inputs
	reg [4:0] opcode;
	reg [31:0] instruction;
	reg bcond;
	reg clk;
	reg rst;

	// Outputs
	wire [4:0]curr_state;
	wire [11:0] micro;
	wire sz_ex;
	wire [31:0] immediate;	
	wire pc_update;
	wire load_ir;
	wire load_mdr;
	wire mem_sel;
	wire mem_wr_en;
	wire reg_file_wr_en;
	wire wr_reg_mux_sel;
	wire op1_sel;
	wire [1:0] op2_sel;
	wire [1:0] alu_demux;
	wire [4:0] alu_ctrl;
	wire [1:0] memory_size;

	// Instantiate the Unit Under Test (UUT)
	cntl_mc uut (
		.instruction(instruction), 
		.bcond(bcond), 
		.clk(clk), 
		.rst(rst), 
		.sz_ex(sz_ex), 
		.immediate(immediate), 
		.mem_sel(mem_sel), 
		.pc_update(pc_update), 
		.load_ir(load_ir), 
		.load_mdr(load_mdr), 
		.mem_wr_en(mem_wr_en), 
		.reg_file_wr_en(reg_file_wr_en), 
		.wr_reg_mux_sel(wr_reg_mux_sel), 
		.op1_sel(op1_sel), 
		.op2_sel(op2_sel), 
		.alu_demux(alu_demux), 
		.alu_ctrl(alu_ctrl), 
		.memory_size(memory_size),
		.curr_state(curr_state),
		.micro(micro)
	);

	initial begin
		// Initialize Inputs
		
		instruction = 0;
		bcond = 0;
		clk = 0;
		rst = 0;

		// Wait 100 ns for global reset to finish
		#2; 
		rst=1;
		#5 rst=0;
		instruction=32'b00000000000000000000000000110100;
		
		#70 $finish;
		
		/*
		instruction=32'b00000000000000000000000000010100;
		instruction=32'b00000000000000000000000001101100;
		instruction=32'b00000000000000000000000001100100;
		instruction=32'b00000000000000000000000001100000;
		instruction=32'b00000000000000000000000000000000;
		instruction=32'b00000000000000000000000000100000;
		instruction=32'b00000000000000000000000000010000;
		instruction=32'b00000000000000000000000000110000;*/

		
        
		// Add stimulus here

	end
      
		always
			#3 clk=~clk;
endmodule
